
typedef uvm_sequencer #(axi4_master_seq_item) axi4_master_seqr;
typedef uvm_sequencer #(axi4_slave_seq_item)  axi4_slave_seqr;
